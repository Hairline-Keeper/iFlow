module Switch_xor(
  input A,
  input B,
  output Y
);
  assign Y =  A ^ B;
endmodule

